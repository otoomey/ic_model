module tb ();

endmodule;
